module rtda

pub struct Slot {
mut:
	num int
	ref &Object
}
