module rtda

struct Slot {
mut:
	num int
	ref &Object
}
