module constant

m
