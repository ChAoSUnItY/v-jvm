module instructions

import vjvm.instructions.constant

__global (
)
