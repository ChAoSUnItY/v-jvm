module instruction

import vjvm.instruction.constant { NOP }

__global (
	nop = &NOP{}
)
