module rtda

pub struct Object {
	// TODO
}
