module vjvm

pub const (
	version = '0.0.1'
)
