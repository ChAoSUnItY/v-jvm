module instructions

import vjvm.instructions.constant
