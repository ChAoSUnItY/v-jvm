module classfile

pub struct ClassFile {
}
