module instructions

import vjvm.instructions.constant { NOP }

__global (
	nop = &NOP{}
)
