module rtda

struct Object {
	// TODO
}
